module testbench();

   tb_full_adder tb0();
      
endmodule
