module alu
  #(parameter xlen = 64)
   ( 
