module uart_tx #(parameter word_size = 8)
   (output serial_out,
    input [word_size-1:0] data_bus,
    input 		  load_xmt_datareg, byte_ready, t_byte, clk, rst_b);


   endmodule
